LIBRARY ieee; 
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

ENTITY OnBoard IS
	PORT (SW		: IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
			KEY	: IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
			LEDR	: OUT	STD_LOGIC_VECTOR(9 DOWNTO 0));
END OnBoard;

ARCHITECTURE Behavior OF OnBoard IS

COMPONENT part1 IS
	PORT (DIN : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			Resetn, Clock, Run : IN STD_LOGIC;
			Done : BUFFER STD_LOGIC;
			BusWires : BUFFER STD_LOGIC_VECTOR(8 DOWNTO 0));
END COMPONENT;

BEGIN

SimpleProcessor : part1 PORT MAP (SW(8 DOWNTO 0), KEY(0), KEY(1), SW(9), LEDR(9), LEDR(8 DOWNTO 0));

END Behavior;