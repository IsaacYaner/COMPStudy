LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part4 IS
	PORT (CLOCK_50	: IN	STD_LOGIC;
			HEX0		: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0));
END part4;

ARCHITECTURE Behavior OF part4 IS

COMPONENT MHZ5 IS
	PORT (CLK	: IN	STD_LOGIC;
			Cout	: OUT	STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT Hnum IS
	PORT (N0					:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			Cin				:	IN		STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

SIGNAL numb : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
	Flash : MHZ5 PORT MAP (CLOCK_50, numb);
	Displ : Hnum PORT MAP (HEX0, numb);
END Behavior;