library verilog;
use verilog.vl_types.all;
entity syncnt8_vlg_vec_tst is
end syncnt8_vlg_vec_tst;
