LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part1 IS
	PORT (HEX0, HEX1	:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			SW				:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0));
END part1;

ARCHITECTURE Behavior OF part1 IS

BEGIN
	HEX0(0)<=(NOT(SW(3)) AND NOT(SW(2)) AND NOT(SW(1)) AND SW(0)) OR (NOT(SW(3)) AND SW(2) AND NOT(SW(1)) AND NOT(SW(0)));
	HEX0(1)<=(NOT(SW(3)) AND SW(2) AND NOT(SW(1)) AND SW(0)) OR (NOT(SW(3)) AND SW(2) AND SW(1) AND NOT(SW(0)));
	HEX0(2)<=(NOT(SW(3)) AND NOT(SW(2)) AND SW(1) AND NOT(SW(0)));
	HEX0(3)<=(NOT(SW(3)) AND NOT(SW(2)) AND NOT(SW(1)) AND SW(0)) OR (NOT(SW(3)) AND SW(2) AND NOT(SW(1)) AND NOT(SW(0))) OR (NOT(SW(3)) AND SW(2) AND SW(1) AND SW(0));
	HEX0(4)<=(NOT(SW(3)) AND SW(0)) OR (NOT(SW(3)) AND SW(2) AND NOT(SW(1)) AND NOT(SW(0))) OR (NOT(SW(2)) AND NOT(SW(1)) AND SW(0));
	HEX0(5)<=(NOT(SW(3)) AND NOT(SW(2)) AND SW(0)) OR (NOT(SW(3)) AND NOT(SW(2)) AND SW(1)) OR (NOT(SW(3)) AND SW(1) AND NOT(SW(0)));
	HEX0(6)<=(NOT(SW(3)) AND NOT(SW(2)) AND NOT(SW(1))) OR (NOT(SW(3)) AND SW(2) AND SW(1) AND SW(0));
END Behavior;