LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part4 IS
	PORT (SW		: IN	STD_LOGIC_VECTOR(8 DOWNTO 0);
			LEDR	: OUT	STD_LOGIC_VECTOR(8 DOWNTO 0);
			LEDG	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			HEX0, HEX1, HEX2, HEX3	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0));
END part4;

ARCHITECTURE Behavior OF part4 IS

COMPONENT Fadder4 IS
	PORT (a, b	: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
			cin	: IN	STD_LOGIC						 ;
			s		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0); 
			cout	: OUT	STD_LOGIC						);
END COMPONENT;

COMPONENT numb IS
	PORT (N0				: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			Cin			: IN		STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT FBCD IS 
	PORT (SW				: IN	STD_LOGIC_VECTOR(4 DOWNTO 0);
			HEX0, HEX1	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			Err			: OUT STD_LOGIC						);
END COMPONENT;
			
SIGNAL Sum : STD_LOGIC_VECTOR(4 DOWNTO 0);
			
--Print the error message
BEGIN
	Disp0 : numb  PORT MAP (HEX3, SW(7 DOWNTO 4));
	Disp1 : numb  PORT MAP (HEX2, SW(3 DOWNTO 0));
	Disp2 : FBCD  PORT MAP (Sum , HEX0, HEX1, LEDG(7));	-- Why could I have larger SW?
	
	Sumup : Fadder4 PORT MAP (SW(7 DOWNTO 4), SW(3 DOWNTO 0), SW(8), Sum(3 DOWNTO 0), Sum(4));
	
END Behavior;