LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part2 IS
	PORT (SW				: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
			HEX0, HEX1	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0));
END part2;

ARCHITECTURE Behavior OF part2 IS

COMPONENT BCDis IS 
	PORT (SW				: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
			HEX0, HEX1	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0));
END COMPONENT;

BEGIN
	Display : BCDis PORT MAP (SW, HEX0, HEX1);
	
END Behavior;