library verilog;
use verilog.vl_types.all;
entity part1q6_vlg_vec_tst is
end part1q6_vlg_vec_tst;
