LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part1 IS
	PORT (HEX0, HEX1	:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			SW				:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0));
END part1;

ARCHITECTURE Behavior OF part1 IS

COMPONENT numb IS	
	PORT (N0					:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			Cin				:	IN		STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

SIGNAL firs, secn : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

firs <= SW(3 DOWNTO 0);
secn <= SW(7 DOWNTO 4);

	Calc0: numb PORT MAP (HEX0, firs);

	Calc1: numb PORT MAP (HEX1, secn);

END Behavior;