LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part3 IS
	PORT (SW		: IN	STD_LOGIC_VECTOR(8 DOWNTO 0);
			LEDR	: OUT	STD_LOGIC_VECTOR(8 DOWNTO 0);
			LEDG	: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END part3;

ARCHITECTURE Behavior OF part3 IS

COMPONENT Fadder4 IS
	PORT (a, b	: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
			cin	: IN	STD_LOGIC						 ;
			s		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0); 
			cout	: OUT	STD_LOGIC						);
END COMPONENT;

BEGIN
	LEDR <= SW;
	AddFour : Fadder4 PORT MAP (SW(7 DOWNTO 4), SW(3 DOWNTO 0), SW(8), LEDG(3 DOWNTO 0), LEDG(4));
	
END Behavior;