library verilog;
use verilog.vl_types.all;
entity divby3_vlg_vec_tst is
end divby3_vlg_vec_tst;
