library verilog;
use verilog.vl_types.all;
entity OnBoard_vlg_vec_tst is
end OnBoard_vlg_vec_tst;
