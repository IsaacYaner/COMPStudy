LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part4 IS
	PORT (SW		: IN	STD_LOGIC_VECTOR(8 DOWNTO 0);
			LEDR	: OUT	STD_LOGIC_VECTOR(8 DOWNTO 0);
			LEDG	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			HEX0, HEX1, HEX2, HEX3	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0));
END part4;

ARCHITECTURE Behavior OF part4 IS

COMPONENT Fadder4 IS
	PORT (a, b	: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
			cin	: IN	STD_LOGIC						 ;
			s		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0); 
			cout	: OUT	STD_LOGIC						);
END COMPONENT;

COMPONENT numb IS
	PORT (N0					:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			Cin				:	IN		STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

BEGIN

END Behavior;